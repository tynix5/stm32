module button(input switch, output led);

assign led = switch;

endmodule